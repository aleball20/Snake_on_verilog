module numbers (number_pixel, clock_25, number_count, selected_number);

/*per permettere la lettura dei numeri, le celle sono di dimensione 10x10 pixel. Quindi ogni quadrato ha 100 bit.
di conseguenza ogni figura Ã¨ rappresentata con 200 bit (2 per ogni pixel). La lettura avviene partendo  
dalla coppie dei 2 MSB che rappresentano il pixel [1][1], per poi procedere leggendo il pixel successivo [2][1]
e cosi via. In uscita si ha un vettore di 2 bit raffigurante il colore del pixel selezionato */
input clock_25;
input [3:0] selected_number;   //Tramite selective decido quale numero prelevare dalla ROM
input [7:0]number_count;              
output number_pixel;
reg [99:0] num[0:15];
reg [99:0] s;

initial begin

    
num[0] = 100'b1111111111100000000110000000011000000001100000000110000000011000000001100000000110000000011111111111; // 0
num[1] = 100'b0000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001; // 1
num[2] = 100'b1111111111000000000100000000010000000001111111111110000000001000000000100000000010000000001111111111; // 2
num[3] = 100'b1111111111000000000100000000010000000001001111111100000000010000000001000000000100000000011111111111; // 3
num[4] = 100'b1000000001100000000110000000011000000001111111111100000000010000000001000000000100000000010000000001; // 4
num[5] = 100'b1111111111100000000010000000001000000000111111111100000000010000000001000000000100000000011111111111; // 5
num[6] = 100'b1111111111100000000010000000001000000000111111111110000000011000000001100000000110000000011111111111; // 6
num[7] = 100'b1111111111000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001; // 7
num[8] = 100'b1111111111100000000110000000011000000001111111111110000000011000000001100000000110000000011111111111; // 8
num[9] = 100'b1111111111100000000110000000011000000001111111111100000000010000000001000000000100000000010000000001; // 9


num[10] = 100'd0;
num[11] = 100'd0;
num[12] = 100'd0;
num[13] = 100'd0;
num[14] = 100'd0;
num[15] = 100'd0;



end


always @ (posedge clock_25)
	begin
			s<= num[selected_number];
	end

assign number_pixel= s[99-number_count];



endmodule