module new_game(clock_25, selected_letter, letter_count);



input clock_25;
input [3:0]selected_letter;
output reg [399:0]letter_count;
reg [399:0] letter[7:0];

initial begin//0 negro y 1 verde usando celdas 20x20 de 1 bit cada una

   
    letter[0]=400'b1111110000000000011111111110000000000111111101110000000001111111001110000000011111100001110000000111111000001110000001111110000001110000011111100000001110000111111000000001110001111110000000001110011111100000000001100111111000000000001001111110000000000001111111100000000000001111111000000000000001111110000000000000011111100000000000000011111000000000000000010000000000000000000000000000000000000000; // N
    letter[1]=400'b1111111111111111111111111111111111111111111000000000000000001110000000000000000011100000000000000000111000000000000000001111111111111110000011111111111111100000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000; // E
    letter[2]=400'b1110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001111110000000000000011111100000011000000111111000001111000001111110000110011000011111100011000011000111111001100000011001111110110000000011011111111000000000001111111000000000000001110000000000000000000000000000000000000000; // W

    letter[3]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // 

    letter[4]=400'b0000001111111111000000011111111111111100001111000000000011100111000000000000001111100000000000000001111000000000000000001110000000000000000011100000000111111110111000000001111111101110000000000000001111100000000000000011011100000000000000110011110000000000011100011111111111111110000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // G
    letter[5]=400'b00000000011100000000 0000000011111000000000000001111111000000000000111001111000000000011100001111000000001110000001111000000111000000001111000011111111111111111001111111111111111111011100000000000001111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000011011000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // A
    letter[6]=400'b1110000000000000011111110000000000001111111110000000000111111110110000000011011111100110000001100111111000110000110001111110000110011000011111100000111100000111111000000110000001111110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // M 
    letter[7]=400'b1111111111111111111111111111111111111111111000000000000000001110000000000000000011100000000000000000111000000000000000001111111111111110000011111111111111100000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000; // E

end


always @ (posedge clock_25)

	begin
		 selected_letter <= letter[selected_letter];
	end



endmodule