/*ROM for printing the name TIME: and SCORE:*/

module rom_background (x_count ,y_count, data, clock_25);
input [7:0] x_count;
input [3:0] y_count;
input clock_25;
output data;
reg [141:0] data_pixel [15:0];
reg [141:0] q;



initial begin
        data_pixel[0] = 142'b111111111111100111100001111110000000011111000011111111110000000001111111100000001111111100000001111111000000011111111110000001111111111000000;
        data_pixel[1] = 142'b111111111111100111100001111110000000111111000011111111110000000111111111100000011111111100000111111111110000011111111111000001111111111000000;
        data_pixel[2] = 142'b111111111111100111100001111111000000111111000011111111110000001111111111100001111111111100001111111111111000011111111111100001111111111000000;
        data_pixel[3] = 142'b000011111000000111100001111111000001111111000011110000000000001111100000000001111110000100011111100011111100011110000111100001111000000000000;
        data_pixel[4] = 142'b000011111000000111100001111111000001111111000011110000000000001111000000000011111000000000011110000001111100011110000111100001111000000000000;
        data_pixel[5] = 142'b000011111000000111100001111111100001111111000011110000000011111111100000000011110000000000111110000000111100011110000111100001111000000001111;
        data_pixel[6] = 142'b000011111000000111100001111111100011111111000011110000000011111111111000000111110000000000111100000000111100011110000111100001111000000001111;
        data_pixel[7] = 142'b000011111000000111100001111011100011101111000011111111100011110111111110000111100000000000111100000000111110011111111111000001111111110001111;
        data_pixel[8] = 142'b000011111000000111100001111011110011101111000011111111100001100011111111000111100000000000111100000000111110011111111110000001111111110000110;
        data_pixel[9] = 142'b000011111000000111100001111011110111101111000011111111100000000000111111100111110000000000111100000000111110011111111110000001111111110000000;
        data_pixel[10] = 142'b000011111000000111100001111001111111001111000011110000000000000000001111110111110000000000111110000000111100011110011111000001111000000000000;
        data_pixel[11] = 142'b000011111000000111100001111001111111001111000011110000000000000000000111110011110000000000111110000000111100011110001111000001111000000000000;
        data_pixel[12] = 142'b000011111000000111100001111000111111001111000011110000000000001000000111110011111100000000011111000011111100011110001111100001111000000000000;
        data_pixel[13] = 142'b000011111000000111100001111000111110001111000011111111100011111111111111100001111111111100001111111111111000011110000111110001111111110001111;
        data_pixel[14] = 142'b000011111000000111100001111000111110001111000011111111110011111111111111100000111111111100000111111111110000011110000011110001111111111001111;
        data_pixel[15] = 142'b000011111000000111100001111000011110001111000011111111110011111111111111000000011111111100000011111111100000011110000011111001111111111001111;
end

always @ (posedge clock_25)
	begin
		q <= data_pixel[y_count];
	end

assign data = q[141-x_count];

endmodule