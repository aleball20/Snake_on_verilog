module game_over(clock_25, selected_letter_over, letter_count_over);



input clock_25;
input [3:0]selected_letter_over;
output reg [399:0]letter_count_over;
reg [399:0] letter_over[15:0];

initial begin//0 negro y 1 verde usando celdas 20x20 de 1 bit cada una

    letter_over[0]=400'b0000001111111111000000011111111111111100001111000000000011100111000000000000001111100000000000000001111000000000000000001110000000000000000011100000000111111110111000000001111111101110000000000000001111100000000000000011011100000000000000110011110000000000011100011111111111111110000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // G
    letter_over[1]=400'b00000000011100000000 0000000011111000000000000001111111000000000000111001111000000000011100001111000000001110000001111000000111000000001111000011111111111111111001111111111111111111011100000000000001111110000000000000001111100000000000000011111000000000000000111110000000000000001111100000000000000011011000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // A
    letter_over[2]=400'b1110000000000000011111110000000000001111111110000000000111111110110000000011011111100110000001100111111000110000110001111110000110011000011111100000111100000111111000000110000001111110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // M 
    letter_over[3]=400'b1111111111111111111111111111111111111111111000000000000000001110000000000000000011100000000000000000111000000000000000001111111111111110000011111111111111100000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000; // E

    letter_over[4]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // 

    letter_over[5]=400'b0000111111111111000000111111111111111000011110000000000111100111000000000000111001110000000000001110011000000000000001100110000000000000011001100000000000000110011000000000000001100110000000000000011001110000000000001110011100000000000011100111000000000000111001110000000000001110011100000000000011100111100000000001111000111111111111111000000011111111111100000000000000000000000000000000000000000000; // O
    letter_over[6]=400'b1110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001111110000000000000011111100000000000000111111000000000000001111110000000000000111001110000000000011100001110000000001110000000111000000111000000000011100011100000000000000111000000000000000000000000000000000000000000000000; // V
    letter_over[7]=400'b1111111111111111111111111111111111111111111000000000000000001110000000000000000011100000000000000000111000000000000000001111111111111110000011111111111111100000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011100000000000000000111000000000000000001110000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000; // E
    letter_over[8]=400'b 111111111111111100001111111111111111100011100000000000001100111000000000000011001110000000000000110011111111111111110000111111111111111110001110000000000000110011100000000000001100111000000000000011001110000000000000110011100000000000001100111000000000000011001110000000000000110011100000000000001100111000000000000011001110000000000000110011100000000000001100000000000000000000000000000000000000000; // R

    letter_over[9]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    letter_over[10]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    letter_over[11]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    letter_over[12]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    letter_over[13]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    letter_over[14]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    letter_over[15]=400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;



end


always @ (posedge clock_25)

	begin
		 selected_letter_over <= letter_over[selected_letter_over];
	end



endmodule