module rom_start_game (x_count ,y_count, data_start_game, clock_25);
input [8:0] x_count;
input [6:0] y_count;
input clock_25;
output data_start_game;
reg [259:0] image_array [65:0];
reg [259:0] q;

initial begin
        image_array[0]  = 260'b00000001010101000000101010101010101010100000000001010100000000000000101010101010000000000101010101010101010100000000000000000000000001010101000000000000000001010100000000000000101010100000000000000010101010000000101010101010100;
        image_array[1]  = 260'b00001111111111110001111111111111111111111000000111111110000000000001111111111111111000001111111111111111111111000000000000000000011111111111111000000000000011111111000000000000111111111000000000000111111111000000111111111111111;
        image_array[2]  = 260'b00111111111111111001111111111111111111110000000111111111000000000001111111111111111100000111111111111111111110000000000000000001111111111111111000000000000111111111000000000001111111111000000000001111111111000000111111111111111;
        image_array[3]  = 260'b01111111111111110001111111111111111111110000000111111111000000000001111111111111111110001111111111111111111111000000000000000011111111111111111000000000000111111111000000000000111111111000000000001111111110000000111111111111111;
        image_array[4]  = 260'b01111111111111111001111111111111111111111000001111111111000000000001111111111111111111000111111111111111111110000000000000000111111111111111111100000000000111111111100000000001111111111100000000001111111111000000111111111111111;
        image_array[5]  = 260'b11111111000001110000000000111111100001000000001111111111100000000001111110000011111111000100001011111100001000000000000000001111111110101011111000000000001111111111100000000000111111111100000000011111111111000000111110000000000;
        image_array[6]  = 260'b11111100000000001000000000111111100000000000011111111111100000000001111110000000111111000000000011111100000000000000000000011111111000000000001000000000001111111111110000000001111111111110000000011111111111000000111110000000000;
        image_array[7]  = 260'b11111100000000000000000000011111100000000000001111011111110000000001111110000001111111000000000111111100000000000000000000011111110000000000000000000000001111101111110000000000111111111100000000011111111110000000111110000000000;
        image_array[8]  = 260'b11111100000000000000000000111111000000000000011111101111100000000001111110000000111111100000000011111100000000000000000000111111100000000000000000000000011111101111110000000001111110111111000000111110111111000000111110000000000;
        image_array[9]  = 260'b11111110000000000000000000011111100000000000111111000111110000000001111110000000111111000000000011111100000000000000000000111111000000000000000000000000011111000111111000000000111110111110000000111111111111000000111110000000000;
        image_array[10] = 260'b11111111100000000000000000111111100000000000111111001111111000000001111110000001111110000000000111111100000000000000000001111111000000000000000000000000111111000111110000000001111110111111000001111100111111000000111110001000000;
        image_array[11] = 260'b11111111111100000000000000011111100000000000111110000111111000000001111111010111111110000000000011111100000000000000000000111111000001010101001000000000111111000111111100000000111110111111000001111101111110000000111111111111110;
        image_array[12] = 260'b01111111111110000000000000111111100000000001111110000111111000000001111111111111111100000000000011111100000000000000000001111110000001111111111110000000111110000011111000000001111110011111100001111100111111000000111111111111110;
        image_array[13] = 260'b00111111111111100000000000011111000000000001111110000011111100000001111111111111111000000000000111111100000000000000000001111111000001111111111100000001111110000111111100000000111110011111100001111001111111000000111111111111110;
        image_array[14] = 260'b00001111111111110000000000111111100000000001111100000111111100000001111111111111100000000000000011111000000000000000000001111110000001111111111110000001111110000011111110000001111110001111100011111000111111000000111111111111110;
        image_array[15] = 260'b00000011111111111000000000011111100000000011111100000011111100000001111111111111110000000000000011111100000000000000000001111111000001111111111110000001111100000001111100000000111110001111110011111001111110000000111111111111110;
        image_array[16] = 260'b00000000111111111000000000111111100000000011111111101011111110000001111110011111110000000000000111111100000000000000000000111111000000001011111100000011111111101111111110000001111110001111100111110000111111000000111110000000000;
        image_array[17] = 260'b00000000001111111100000000011111100000000111111111111111111110000001111110000111111100000000000011111100000000000000000001111111000000000011111110000011111111111111111111000000111110001111111011110001111111000000111111000000000;
        image_array[18] = 260'b00000000000111111100000000111111000000000111111111111111111110000001111110000111111100000000000011111100000000000000000000111111100000000001111100000111111111111111111110000001111110000111111111110000111111000000111110000000000;
        image_array[19] = 260'b00000000000111111100000000011111100000000111111111111111111111000001111110000011111110000000000111111100000000000000000000111111100000000011111110000111111111111111111111000000111110000111111111100001111110000000111111000000000;
        image_array[20] = 260'b10000000000111111100000000111111100000001111111111111111111111000001111110000001111111000000000011111100000000000000000000011111111000000011111100000111111111111111111111100001111110000011111111100000111111000000111110000000000;
        image_array[21] = 260'b01110000001011111100000000001111110000000111111000000000011111100000111111000000111111100000000001111110000000000000000000001111111111010101111111000111111100000000011111110000011111000001111111110000111111100000111111100000000;
        image_array[22] = 260'b01111111111111111100000000011111100000000111111000000000011111110000111111000000011111110000000011111110000000000000000000000111111111111111111111000111111000000000001111110000111111000001111111100000011111100000111111111111111;
        image_array[23] = 260'b01111111111111111000000000001111110000001111111000000000001111110000111111000000001111110000000001111110000000000000000000000011111111111111111110000111111000000000001111110000011111000000111111100000111111000000111111111111111;
        image_array[24] = 260'b01111111111111111000000000011111110000001111110000000000001111111000111111000000001111111000000011111100000000000000000000000001111111111111111111001111111000000000001111111000111111000000111111000000011111100000111111111111111;
        image_array[25] = 260'b01111111111111100000000000001111110000011111110000000000001111110000111111000000001111111100000001111110000000000000000000000000011111111111111000001111110000000000000111111000011111000000011111100000111111100000111111111111111;
        image_array[26] = 260'b00010111110100000000000000001101100000001011010000000000000111011000101101000000000011011000000001101100000000000000000000000000000010111101000000001011010000000000000110111000111011000000110110000000010111000000111111111111111;
        image_array[27] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[28] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[29] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[30] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[31] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[32] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[33] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[34] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[35] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[36] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[37] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[38] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[39] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[40] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[41] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[42] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[43] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[44] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[45] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[46] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[47] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[48] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[49] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[50] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[51] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[52] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[53] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[54] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[55] = 260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        image_array[56] = 260'b00000000000000000000000000000000000000000000000000000000000000010110110101011011010101101101011011010011011010000000010100001010001010101000101000010100011011011011011000010100000000000000000000000000000000000000000000000000000;
        image_array[57] = 260'b00000000000000000000000000000000000000000000000000000000000000011111111101111111110111111111111111110111111110000000111110001111011111111001111000011101011111111111111100111100000000000000000000000000000000000000000000000000000;
        image_array[58] = 260'b00000000000000000000000000000000000000000000000000000000000000011110111111111011110111101011111010101111010100000000111110001111001111111001110000011110111011110101011100111000000000000000000000000000000000000000000000000000000;
        image_array[59] = 260'b00000000000000000000000000000000000000000000000000000000000000001110001110110001111111000001111000000111000000000001111111001111111110111011110000011101111011101000011110111000000000000000000000000000000000000000000000000000000;
        image_array[60] = 260'b00000000000000000000000000000000000000000000000000000000000000011110011111111001110111111100111111101111111101000001110111001111101110011111100000011111110011111110001111110000000000000000000000000000000000000000000000000000000;
        image_array[61] = 260'b00000000000000000000000000000000000000000000000000000000000000011111011101111111111111111101111111110111111110000001110111011111111110011111000000011111110011111111000111110000000000000000000000000000000000000000000000000000000;
        image_array[62] = 260'b00000000000000000000000000000000000000000000000000000000000000011111111110111111100111001000000101111000101111000011111111101110111110001111000000011111110011100000000111100000000000000000000000000000000000000000000000000000000;
        image_array[63] = 260'b00000000000000000000000000000000000000000000000000000000000000001110000001111011110111100100010001110010001111000011111111101110111110001111000000011101111011110101000111100000000000000000000000000000000000000000000000000000000;
        image_array[64] = 260'b00000000000000000000000000000000000000000000000000000000000000011100010001110011110111111111111111111111111110000011100111111110011111000110000000011100111111111111000011100000000000000000000000000000000000000000000000000000000;
        image_array[65] = 260'b00000000000000000000000000000000000000000000000000000000000000011110000001111001101011111110111111101011111110000111100001110110011110001111000000011100111011111111100011000000000000000000000000000000000000000000000000000000000;
end

always @ (posedge clock_25)
	begin
		q <= image_array[y_count];
	end

assign data_start_game = q[259-x_count];

endmodule