module rom_game_over (x_count ,y_count, data_game_over, clock_25);
input [7:0] x_count;
input [4:0] y_count;
input clock_25;
output data_game_over;
reg [183:0] image_array [22:0];
reg [183:0] q;



initial begin
    
        image_array[0] =  184'b0000000001111110100000000000001111110000000000011111100000000000011111110000001111111111110000000000000000000011111010000000011111000000000001111000011111111111100000111111111101000000;
        image_array[1] =  184'b0000001111111111111000000000011111110000000000111111111000000000111111110000011111111111110000000000000000011111111111000000001111100000000011111100011111111111110000111111111111100000;
        image_array[2] =  184'b0000111111111111111000000000011111111000000000011111111000000000111111110000011111111111110000000000000000111111111111110000011111100000000011111000011111111111110001111111111111111000;
        image_array[3] =  184'b0001011111111111111000000000011111111000000000111111111000000000111111111000001111111111111000000000000001111111111111111000001111100000000011111000011111111111110000111111011111111000;
        image_array[4] =  184'b0001111111100101111000000000111111111000000000011111111000000001111111110000011111010010010000000000000011111111011111111100001111110000000111111000011111001001000000111110000111111100;
        image_array[5] =  184'b0011111100000000001000000000111101111100000000111111111100000001111111110000011111000000000000000000000111111100000011111100000111110000000111110000011111000000000001111110000011111100;
        image_array[6] =  184'b0011111101000000000000000001111111111000000000111111111000000011101111110000111111000000000000000000001111110000000011111100001111100000001111100000111110000000000001111100000011111000;
        image_array[7] =  184'b0111111000000000000000000001111100111110000000111110111110000011111111110000001111000000000000000000001111110000000001111110000111111000000111110000011111000000000000111110000011111100;
        image_array[8] =  184'b0111111000000000000000000001111100111110000000011110111110000011110111110000011111000000000000000000001111110000000000111111000011111000001111100000011111000000000001111110000001111000;
        image_array[9] =  184'b1111110000000000000000000011110001111100000001111101111100000111101111110000111111000000000000000000011111000000000001111110000111110000011111000000111110000000000001111100000111111000;
        image_array[10] = 184'b1111100000010101010100000011111000111110000000011110011111000111100111110000011111111111110000000000001111100000000000111111000011111100001111100000011111111111110000111110010111111000;
        image_array[11] = 184'b1111110000111111111100000011111000011111000000111110011110000111110111110000001111111111110000000000001111100000000000011110000001111000011111000000011111111111100001111111111111110000;
        image_array[12] = 184'b1111100000111111111100000111110000011111000000011110011111000111100111111000011111111111110000000000011111100000000000111111000001111100011111000000011111111111110000111111111111000000;
        image_array[13] = 184'b1111100000111111111100000111110000011111100000111110001111101111000111110000011111111111100000000000001111100000000000111111000001111110011111000000011111111111100000111111111111000000;
        image_array[14] = 184'b1111110000010111111100000111111010111111100000011110011111101111100111110000011111000000000000000000001111110000000000111110000000111100111110000000011111000000000000111110111111100000;
        image_array[15] = 184'b0111110000000001111100000111111111111111100000111110000111101111000111111000001111000000000000000000001111110000000000111111000000111110111110000000011111000000000001111110001111110000;
        image_array[16] = 184'b1111111000000011111100001111111111111111110000011110001111111110000111110000011111100000000000000000001111110000000001111110000000111110111110000000011111000000000000111110001111110000;
        image_array[17] = 184'b0111111000000001111100001111111111111111110000111110000111111110000111110000011111000000000000000000000111111000000011111100000000111111111100000000011111000000000000111110000111111000;
        image_array[18] = 184'b0011111110100011111100011111101010101111110000011110000111111110000111111000011111100000000000000000000111111110010111111100000000011111111100000000011111000000000000111110000011111100;
        image_array[19] = 184'b0011111111111111111100011111100000000111111000111110000011111100000111110000001111111111111000000000000011111111111111111000000000011111111100000000011111111111110001111110000001111100;
        image_array[20] = 184'b0001111111111111111100011111000000000011111000011110000011111110000111110000011111111111111000000000000001111111111111110000000000001111111000000000011111111111110000111110000001111110;
        image_array[21] = 184'b0000111111111111111100111111000000000011111000111110000011111100000111111000011111111111111000000000000000111111111111010000000000001111111000000000011111111111110000111110000001111110;
        image_array[22] = 184'b0000000111111111100000111111000000000011111100011110000001111000000111110000011111111111111000000000000000001111111101000000000000001111110000000000011111111111111001111110000000111111;   
end

always @ (posedge clock_25)
	begin
		q <= image_array[y_count];
	end

assign data_game_over = q[183-x_count];

endmodule